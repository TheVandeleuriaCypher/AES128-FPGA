`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Engineer: Jason Li
// 
// Module Name:  InvMixColumns
// Project Name: AES128
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//Step 1) Takes input of an 128 bit number, inData
//Step 2) Performs matrix multiplication with the inverse matrix counterpart to MixColumns
//Step 3) Calls the mult functio when the matrices are expanded, as we need to account for 
//Step 4) Returns it as outData
//////////////////////////////////////////////////////////////////////////////////
module InvMixColumns(
	 input [127:0] inData,
	 output [127:0] outData
    );
	 
	 wire [7:0] s0,s1,s2,s3,s4,s5,s6,s7,s8,s9,s10,s11,s12,s13,s14,s15;
	 reg [7:0] t0,t1,t2,t3,t4,t5,t6,t7,t8,t9,t10,t11,t12,t13,t14,t15;
	 
	 //assigning variables to inputs
	 assign s0 = inData[7:0];
	 assign s1 = inData[15:8];
	 assign s2 = inData[23:16];
	 assign s3 = inData[31:24];
	 assign s4 = inData[39:32];
	 assign s5 = inData[47:40];
	 assign s6 = inData[55:48];
	 assign s7 = inData[63:56];
	 assign s8 = inData[71:64];
	 assign s9 = inData[79:72];
	 assign s10 = inData[87:80];
	 assign s11 = inData[95:88];
	 assign s12 = inData[103:96];
	 assign s13 = inData[111:104];
	 assign s14 = inData[119:112];
	 assign s15 = inData[127:120];
	 
	 
	 //Step 2
	 //Performs matrix multiplication with the inverse matrix counterpart to MixColumns
	 always @(*)
	 begin
		  t15 = decmult(s15,14) ^ decmult(s14,11) ^ decmult(s13,13) ^ decmult(s12,9);
		  t14 = decmult(s15,9) ^ decmult(s14,14) ^ decmult(s13,11) ^ decmult(s12,13);
		  t13 = decmult(s15,13) ^ decmult(s14,9) ^ decmult(s13,14) ^ decmult(s12,11);
		  t12 = decmult(s15,11) ^ decmult(s14,13) ^ decmult(s13,9) ^ decmult(s12,14);
		  
		  t11 = decmult(s11,14) ^ decmult(s10,11) ^ decmult(s9,13) ^ decmult(s8,9);
		  t10 = decmult(s11,9) ^ decmult(s10,14) ^ decmult(s9,11) ^ decmult(s8,13);
		  t9 = decmult(s11,13) ^ decmult(s10,9) ^ decmult(s9,14) ^ decmult(s8,11);
		  t8 = decmult(s11,11) ^ decmult(s10,13) ^ decmult(s9,9) ^ decmult(s8,14);
		  
		  t7 = decmult(s7,14) ^ decmult(s6,11) ^ decmult(s5,13) ^ decmult(s4,9);
		  t6 = decmult(s7,9) ^ decmult(s6,14) ^ decmult(s5,11) ^ decmult(s4,13);
		  t5 = decmult(s7,13) ^ decmult(s6,9) ^ decmult(s5,14) ^ decmult(s4,11);
		  t4 = decmult(s7,11) ^ decmult(s6,13) ^ decmult(s5,9) ^ decmult(s4,14);
		  
		  t3 = decmult(s3,14) ^ decmult(s2,11) ^ decmult(s1,13) ^ decmult(s0,9);
		  t2 = decmult(s3,9) ^ decmult(s2,14) ^ decmult(s1,11) ^ decmult(s0,13);
		  t1 = decmult(s3,13) ^ decmult(s2,9) ^ decmult(s1,14) ^ decmult(s0,11);
		  t0 = decmult(s3,11) ^ decmult(s2,13) ^ decmult(s1,9) ^ decmult(s0,14);
	 end
	 
	 //assigns the individual t variables to the output variable
	 assign outData[7:0] = t0;
	 assign outData[15:8] = t1;
	 assign outData[23:16] = t2;
	 assign outData[31:24] = t3;
	 assign outData[39:32] = t4;
	 assign outData[47:40] = t5;
	 assign outData[55:48] = t6;
	 assign outData[63:56] = t7;
	 assign outData[71:64] = t8;
	 assign outData[79:72] = t9;
	 assign outData[87:80] = t10;
	 assign outData[95:88] = t11;
	 assign outData[103:96] = t12;
	 assign outData[111:104] = t13;
	 assign outData[119:112] = t14;
	 assign outData[127:120] = t15;
	 
	 //we utilise long case statements in functions to perform the matrix multiplications as the calculations would take signifcantly more calculations
	 function [7:0] decmult(input[7:0] num1,num2);
		  case(num2)
				8'h09: decmult=decmult_9(num1);
				8'h0b: decmult=decmult_11(num1);
				8'h0d: decmult=decmult_13(num1);
				8'h0e: decmult=decmult_14(num1);
		  endcase
	 endfunction
	 
	 //function holding case statement multiply by 9
	 function [7:0] decmult_9(input [7:0] num);
		  case (num)
				8'h00: decmult_9 = 8'h00;
				8'h01: decmult_9 = 8'h09;
				8'h02: decmult_9 = 8'h12;
				8'h03: decmult_9 = 8'h1B;
				8'h04: decmult_9 = 8'h24;
				8'h05: decmult_9 = 8'h2D;
				8'h06: decmult_9 = 8'h36;
				8'h07: decmult_9 = 8'h3F;
				8'h08: decmult_9 = 8'h48;
				8'h09: decmult_9 = 8'h41;
				8'h0A: decmult_9 = 8'h5A;
				8'h0B: decmult_9 = 8'h53;
				8'h0C: decmult_9 = 8'h6C;
				8'h0D: decmult_9 = 8'h65;
				8'h0E: decmult_9 = 8'h7E;
				8'h0F: decmult_9 = 8'h77;
				8'h10: decmult_9 = 8'h90;
				8'h11: decmult_9 = 8'h99;
				8'h12: decmult_9 = 8'h82;
				8'h13: decmult_9 = 8'h8B;
				8'h14: decmult_9 = 8'hB4;
				8'h15: decmult_9 = 8'hBD;
				8'h16: decmult_9 = 8'hA6;
				8'h17: decmult_9 = 8'hAF;
				8'h18: decmult_9 = 8'hD8;
				8'h19: decmult_9 = 8'hD1;
				8'h1A: decmult_9 = 8'hCA;
				8'h1B: decmult_9 = 8'hC3;
				8'h1C: decmult_9 = 8'hFC;
				8'h1D: decmult_9 = 8'hF5;
				8'h1E: decmult_9 = 8'hEE;
				8'h1F: decmult_9 = 8'hE7;
				8'h20: decmult_9 = 8'h3B;
				8'h21: decmult_9 = 8'h32;
				8'h22: decmult_9 = 8'h29;
				8'h23: decmult_9 = 8'h20;
				8'h24: decmult_9 = 8'h1F;
				8'h25: decmult_9 = 8'h16;
				8'h26: decmult_9 = 8'h0D;
				8'h27: decmult_9 = 8'h04;
				8'h28: decmult_9 = 8'h73;
				8'h29: decmult_9 = 8'h7A;
				8'h2A: decmult_9 = 8'h61;
				8'h2B: decmult_9 = 8'h68;
				8'h2C: decmult_9 = 8'h57;
				8'h2D: decmult_9 = 8'h5E;
				8'h2E: decmult_9 = 8'h45;
				8'h2F: decmult_9 = 8'h4C;
				8'h30: decmult_9 = 8'hAB;
				8'h31: decmult_9 = 8'hA2;
				8'h32: decmult_9 = 8'hB9;
				8'h33: decmult_9 = 8'hB0;
				8'h34: decmult_9 = 8'h8F;
				8'h35: decmult_9 = 8'h86;
				8'h36: decmult_9 = 8'h9D;
				8'h37: decmult_9 = 8'h94;
				8'h38: decmult_9 = 8'hE3;
				8'h39: decmult_9 = 8'hEA;
				8'h3A: decmult_9 = 8'hF1;
				8'h3B: decmult_9 = 8'hF8;
				8'h3C: decmult_9 = 8'hC7;
				8'h3D: decmult_9 = 8'hCE;
				8'h3E: decmult_9 = 8'hD5;
				8'h3F: decmult_9 = 8'hDC;
				8'h40: decmult_9 = 8'h76;
				8'h41: decmult_9 = 8'h7F;
				8'h42: decmult_9 = 8'h64;
				8'h43: decmult_9 = 8'h6D;
				8'h44: decmult_9 = 8'h52;
				8'h45: decmult_9 = 8'h5B;
				8'h46: decmult_9 = 8'h40;
				8'h47: decmult_9 = 8'h49;
				8'h48: decmult_9 = 8'h3E;
				8'h49: decmult_9 = 8'h37;
				8'h4A: decmult_9 = 8'h2C;
				8'h4B: decmult_9 = 8'h25;
				8'h4C: decmult_9 = 8'h1A;
				8'h4D: decmult_9 = 8'h13;
				8'h4E: decmult_9 = 8'h08;
				8'h4F: decmult_9 = 8'h01;
				8'h50: decmult_9 = 8'hE6;
				8'h51: decmult_9 = 8'hEF;
				8'h52: decmult_9 = 8'hF4;
				8'h53: decmult_9 = 8'hFD;
				8'h54: decmult_9 = 8'hC2;
				8'h55: decmult_9 = 8'hCB;
				8'h56: decmult_9 = 8'hD0;
				8'h57: decmult_9 = 8'hD9;
				8'h58: decmult_9 = 8'hAE;
				8'h59: decmult_9 = 8'hA7;
				8'h5A: decmult_9 = 8'hBC;
				8'h5B: decmult_9 = 8'hB5;
				8'h5C: decmult_9 = 8'h8A;
				8'h5D: decmult_9 = 8'h83;
				8'h5E: decmult_9 = 8'h98;
				8'h5F: decmult_9 = 8'h91;
				8'h60: decmult_9 = 8'h4D;
				8'h61: decmult_9 = 8'h44;
				8'h62: decmult_9 = 8'h5F;
				8'h63: decmult_9 = 8'h56;
				8'h64: decmult_9 = 8'h69;
				8'h65: decmult_9 = 8'h60;
				8'h66: decmult_9 = 8'h7B;
				8'h67: decmult_9 = 8'h72;
				8'h68: decmult_9 = 8'h05;
				8'h69: decmult_9 = 8'h0C;
				8'h6A: decmult_9 = 8'h17;
				8'h6B: decmult_9 = 8'h1E;
				8'h6C: decmult_9 = 8'h21;
				8'h6D: decmult_9 = 8'h28;
				8'h6E: decmult_9 = 8'h33;
				8'h6F: decmult_9 = 8'h3A;
				8'h70: decmult_9 = 8'hDD;
				8'h71: decmult_9 = 8'hD4;
				8'h72: decmult_9 = 8'hCF;
				8'h73: decmult_9 = 8'hC6;
				8'h74: decmult_9 = 8'hF9;
				8'h75: decmult_9 = 8'hF0;
				8'h76: decmult_9 = 8'hEB;
				8'h77: decmult_9 = 8'hE2;
				8'h78: decmult_9 = 8'h95;
				8'h79: decmult_9 = 8'h9C;
				8'h7A: decmult_9 = 8'h87;
				8'h7B: decmult_9 = 8'h8E;
				8'h7C: decmult_9 = 8'hB1;
				8'h7D: decmult_9 = 8'hB8;
				8'h7E: decmult_9 = 8'hA3;
				8'h7F: decmult_9 = 8'hAA;
				8'h80: decmult_9 = 8'hEC;
				8'h81: decmult_9 = 8'hE5;
				8'h82: decmult_9 = 8'hFE;
				8'h83: decmult_9 = 8'hF7;
				8'h84: decmult_9 = 8'hC8;
				8'h85: decmult_9 = 8'hC1;
				8'h86: decmult_9 = 8'hDA;
				8'h87: decmult_9 = 8'hD3;
				8'h88: decmult_9 = 8'hA4;
				8'h89: decmult_9 = 8'hAD;
				8'h8A: decmult_9 = 8'hB6;
				8'h8B: decmult_9 = 8'hBF;
				8'h8C: decmult_9 = 8'h80;
				8'h8D: decmult_9 = 8'h89;
				8'h8E: decmult_9 = 8'h92;
				8'h8F: decmult_9 = 8'h9B;
				8'h90: decmult_9 = 8'h7C;
				8'h91: decmult_9 = 8'h75;
				8'h92: decmult_9 = 8'h6E;
				8'h93: decmult_9 = 8'h67;
				8'h94: decmult_9 = 8'h58;
				8'h95: decmult_9 = 8'h51;
				8'h96: decmult_9 = 8'h4A;
				8'h97: decmult_9 = 8'h43;
				8'h98: decmult_9 = 8'h34;
				8'h99: decmult_9 = 8'h3D;
				8'h9A: decmult_9 = 8'h26;
				8'h9B: decmult_9 = 8'h2F;
				8'h9C: decmult_9 = 8'h10;
				8'h9D: decmult_9 = 8'h19;
				8'h9E: decmult_9 = 8'h02;
				8'h9F: decmult_9 = 8'h0B;
				8'hA0: decmult_9 = 8'hD7;
				8'hA1: decmult_9 = 8'hDE;
				8'hA2: decmult_9 = 8'hC5;
				8'hA3: decmult_9 = 8'hCC;
				8'hA4: decmult_9 = 8'hF3;
				8'hA5: decmult_9 = 8'hFA;
				8'hA6: decmult_9 = 8'hE1;
				8'hA7: decmult_9 = 8'hE8;
				8'hA8: decmult_9 = 8'h9F;
				8'hA9: decmult_9 = 8'h96;
				8'hAA: decmult_9 = 8'h8D;
				8'hAB: decmult_9 = 8'h84;
				8'hAC: decmult_9 = 8'hBB;
				8'hAD: decmult_9 = 8'hB2;
				8'hAE: decmult_9 = 8'hA9;
				8'hAF: decmult_9 = 8'hA0;
				8'hB0: decmult_9 = 8'h47;
				8'hB1: decmult_9 = 8'h4E;
				8'hB2: decmult_9 = 8'h55;
				8'hB3: decmult_9 = 8'h5C;
				8'hB4: decmult_9 = 8'h63;
				8'hB5: decmult_9 = 8'h6A;
				8'hB6: decmult_9 = 8'h71;
				8'hB7: decmult_9 = 8'h78;
				8'hB8: decmult_9 = 8'h0F;
				8'hB9: decmult_9 = 8'h06;
				8'hBA: decmult_9 = 8'h1D;
				8'hBB: decmult_9 = 8'h14;
				8'hBC: decmult_9 = 8'h2B;
				8'hBD: decmult_9 = 8'h22;
				8'hBE: decmult_9 = 8'h39;
				8'hBF: decmult_9 = 8'h30;
				8'hC0: decmult_9 = 8'h9A;
				8'hC1: decmult_9 = 8'h93;
				8'hC2: decmult_9 = 8'h88;
				8'hC3: decmult_9 = 8'h81;
				8'hC4: decmult_9 = 8'hBE;
				8'hC5: decmult_9 = 8'hB7;
				8'hC6: decmult_9 = 8'hAC;
				8'hC7: decmult_9 = 8'hA5;
				8'hC8: decmult_9 = 8'hD2;
				8'hC9: decmult_9 = 8'hDB;
				8'hCA: decmult_9 = 8'hC0;
				8'hCB: decmult_9 = 8'hC9;
				8'hCC: decmult_9 = 8'hF6;
				8'hCD: decmult_9 = 8'hFF;
				8'hCE: decmult_9 = 8'hE4;
				8'hCF: decmult_9 = 8'hED;
				8'hD0: decmult_9 = 8'h0A;
				8'hD1: decmult_9 = 8'h03;
				8'hD2: decmult_9 = 8'h18;
				8'hD3: decmult_9 = 8'h11;
				8'hD4: decmult_9 = 8'h2E;
				8'hD5: decmult_9 = 8'h27;
				8'hD6: decmult_9 = 8'h3C;
				8'hD7: decmult_9 = 8'h35;
				8'hD8: decmult_9 = 8'h42;
				8'hD9: decmult_9 = 8'h4B;
				8'hDA: decmult_9 = 8'h50;
				8'hDB: decmult_9 = 8'h59;
				8'hDC: decmult_9 = 8'h66;
				8'hDD: decmult_9 = 8'h6F;
				8'hDE: decmult_9 = 8'h74;
				8'hDF: decmult_9 = 8'h7D;
				8'hE0: decmult_9 = 8'hA1;
				8'hE1: decmult_9 = 8'hA8;
				8'hE2: decmult_9 = 8'hB3;
				8'hE3: decmult_9 = 8'hBA;
				8'hE4: decmult_9 = 8'h85;
				8'hE5: decmult_9 = 8'h8C;
				8'hE6: decmult_9 = 8'h97;
				8'hE7: decmult_9 = 8'h9E;
				8'hE8: decmult_9 = 8'hE9;
				8'hE9: decmult_9 = 8'hE0;
				8'hEA: decmult_9 = 8'hFB;
				8'hEB: decmult_9 = 8'hF2;
				8'hEC: decmult_9 = 8'hCD;
				8'hED: decmult_9 = 8'hC4;
				8'hEE: decmult_9 = 8'hDF;
				8'hEF: decmult_9 = 8'hD6;
				8'hF0: decmult_9 = 8'h31;
				8'hF1: decmult_9 = 8'h38;
				8'hF2: decmult_9 = 8'h23;
				8'hF3: decmult_9 = 8'h2A;
				8'hF4: decmult_9 = 8'h15;
				8'hF5: decmult_9 = 8'h1C;
				8'hF6: decmult_9 = 8'h07;
				8'hF7: decmult_9 = 8'h0E;
				8'hF8: decmult_9 = 8'h79;
				8'hF9: decmult_9 = 8'h70;
				8'hFA: decmult_9 = 8'h6B;
				8'hFB: decmult_9 = 8'h62;
				8'hFC: decmult_9 = 8'h5D;
				8'hFD: decmult_9 = 8'h54;
				8'hFE: decmult_9 = 8'h4F;
				8'hFF: decmult_9 = 8'h46;
		  endcase
	 endfunction
	 
	 //function holding case statement multiply by 11
	 function [7:0] decmult_11(input [7:0] num);
		  case (num)
				8'h00: decmult_11 = 8'h00;
				8'h01: decmult_11 = 8'h0B;
				8'h02: decmult_11 = 8'h16;
				8'h03: decmult_11 = 8'h1D;
				8'h04: decmult_11 = 8'h2C;
				8'h05: decmult_11 = 8'h27;
				8'h06: decmult_11 = 8'h3A;
				8'h07: decmult_11 = 8'h31;
				8'h08: decmult_11 = 8'h58;
				8'h09: decmult_11 = 8'h53;
				8'h0A: decmult_11 = 8'h4E;
				8'h0B: decmult_11 = 8'h45;
				8'h0C: decmult_11 = 8'h74;
				8'h0D: decmult_11 = 8'h7F;
				8'h0E: decmult_11 = 8'h62;
				8'h0F: decmult_11 = 8'h69;
				8'h10: decmult_11 = 8'hB0;
				8'h11: decmult_11 = 8'hBB;
				8'h12: decmult_11 = 8'hA6;
				8'h13: decmult_11 = 8'hAD;
				8'h14: decmult_11 = 8'h9C;
				8'h15: decmult_11 = 8'h97;
				8'h16: decmult_11 = 8'h8A;
				8'h17: decmult_11 = 8'h81;
				8'h18: decmult_11 = 8'hE8;
				8'h19: decmult_11 = 8'hE3;
				8'h1A: decmult_11 = 8'hFE;
				8'h1B: decmult_11 = 8'hF5;
				8'h1C: decmult_11 = 8'hC4;
				8'h1D: decmult_11 = 8'hCF;
				8'h1E: decmult_11 = 8'hD2;
				8'h1F: decmult_11 = 8'hD9;
				8'h20: decmult_11 = 8'h7B;
				8'h21: decmult_11 = 8'h70;
				8'h22: decmult_11 = 8'h6D;
				8'h23: decmult_11 = 8'h66;
				8'h24: decmult_11 = 8'h57;
				8'h25: decmult_11 = 8'h5C;
				8'h26: decmult_11 = 8'h41;
				8'h27: decmult_11 = 8'h4A;
				8'h28: decmult_11 = 8'h23;
				8'h29: decmult_11 = 8'h28;
				8'h2A: decmult_11 = 8'h35;
				8'h2B: decmult_11 = 8'h3E;
				8'h2C: decmult_11 = 8'h0F;
				8'h2D: decmult_11 = 8'h04;
				8'h2E: decmult_11 = 8'h19;
				8'h2F: decmult_11 = 8'h12;
				8'h30: decmult_11 = 8'hCB;
				8'h31: decmult_11 = 8'hC0;
				8'h32: decmult_11 = 8'hDD;
				8'h33: decmult_11 = 8'hD6;
				8'h34: decmult_11 = 8'hE7;
				8'h35: decmult_11 = 8'hEC;
				8'h36: decmult_11 = 8'hF1;
				8'h37: decmult_11 = 8'hFA;
				8'h38: decmult_11 = 8'h93;
				8'h39: decmult_11 = 8'h98;
				8'h3A: decmult_11 = 8'h85;
				8'h3B: decmult_11 = 8'h8E;
				8'h3C: decmult_11 = 8'hBF;
				8'h3D: decmult_11 = 8'hB4;
				8'h3E: decmult_11 = 8'hA9;
				8'h3F: decmult_11 = 8'hA2;
				8'h40: decmult_11 = 8'hF6;
				8'h41: decmult_11 = 8'hFD;
				8'h42: decmult_11 = 8'hE0;
				8'h43: decmult_11 = 8'hEB;
				8'h44: decmult_11 = 8'hDA;
				8'h45: decmult_11 = 8'hD1;
				8'h46: decmult_11 = 8'hCC;
				8'h47: decmult_11 = 8'hC7;
				8'h48: decmult_11 = 8'hAE;
				8'h49: decmult_11 = 8'hA5;
				8'h4A: decmult_11 = 8'hB8;
				8'h4B: decmult_11 = 8'hB3;
				8'h4C: decmult_11 = 8'h82;
				8'h4D: decmult_11 = 8'h89;
				8'h4E: decmult_11 = 8'h94;
				8'h4F: decmult_11 = 8'h9F;
				8'h50: decmult_11 = 8'h46;
				8'h51: decmult_11 = 8'h4D;
				8'h52: decmult_11 = 8'h50;
				8'h53: decmult_11 = 8'h5B;
				8'h54: decmult_11 = 8'h6A;
				8'h55: decmult_11 = 8'h61;
				8'h56: decmult_11 = 8'h7C;
				8'h57: decmult_11 = 8'h77;
				8'h58: decmult_11 = 8'h1E;
				8'h59: decmult_11 = 8'h15;
				8'h5A: decmult_11 = 8'h08;
				8'h5B: decmult_11 = 8'h03;
				8'h5C: decmult_11 = 8'h32;
				8'h5D: decmult_11 = 8'h39;
				8'h5E: decmult_11 = 8'h24;
				8'h5F: decmult_11 = 8'h2F;
				8'h60: decmult_11 = 8'h8D;
				8'h61: decmult_11 = 8'h86;
				8'h62: decmult_11 = 8'h9B;
				8'h63: decmult_11 = 8'h90;
				8'h64: decmult_11 = 8'hA1;
				8'h65: decmult_11 = 8'hAA;
				8'h66: decmult_11 = 8'hB7;
				8'h67: decmult_11 = 8'hBC;
				8'h68: decmult_11 = 8'hD5;
				8'h69: decmult_11 = 8'hDE;
				8'h6A: decmult_11 = 8'hC3;
				8'h6B: decmult_11 = 8'hC8;
				8'h6C: decmult_11 = 8'hF9;
				8'h6D: decmult_11 = 8'hF2;
				8'h6E: decmult_11 = 8'hEF;
				8'h6F: decmult_11 = 8'hE4;
				8'h70: decmult_11 = 8'h3D;
				8'h71: decmult_11 = 8'h36;
				8'h72: decmult_11 = 8'h2B;
				8'h73: decmult_11 = 8'h20;
				8'h74: decmult_11 = 8'h11;
				8'h75: decmult_11 = 8'h1A;
				8'h76: decmult_11 = 8'h07;
				8'h77: decmult_11 = 8'h0C;
				8'h78: decmult_11 = 8'h65;
				8'h79: decmult_11 = 8'h6E;
				8'h7A: decmult_11 = 8'h73;
				8'h7B: decmult_11 = 8'h78;
				8'h7C: decmult_11 = 8'h49;
				8'h7D: decmult_11 = 8'h42;
				8'h7E: decmult_11 = 8'h5F;
				8'h7F: decmult_11 = 8'h54;
				8'h80: decmult_11 = 8'hF7;
				8'h81: decmult_11 = 8'hFC;
				8'h82: decmult_11 = 8'hE1;
				8'h83: decmult_11 = 8'hEA;
				8'h84: decmult_11 = 8'hDB;
				8'h85: decmult_11 = 8'hD0;
				8'h86: decmult_11 = 8'hCD;
				8'h87: decmult_11 = 8'hC6;
				8'h88: decmult_11 = 8'hAF;
				8'h89: decmult_11 = 8'hA4;
				8'h8A: decmult_11 = 8'hB9;
				8'h8B: decmult_11 = 8'hB2;
				8'h8C: decmult_11 = 8'h83;
				8'h8D: decmult_11 = 8'h88;
				8'h8E: decmult_11 = 8'h95;
				8'h8F: decmult_11 = 8'h9E;
				8'h90: decmult_11 = 8'h47;
				8'h91: decmult_11 = 8'h4C;
				8'h92: decmult_11 = 8'h51;
				8'h93: decmult_11 = 8'h5A;
				8'h94: decmult_11 = 8'h6B;
				8'h95: decmult_11 = 8'h60;
				8'h96: decmult_11 = 8'h7D;
				8'h97: decmult_11 = 8'h76;
				8'h98: decmult_11 = 8'h1F;
				8'h99: decmult_11 = 8'h14;
				8'h9A: decmult_11 = 8'h09;
				8'h9B: decmult_11 = 8'h02;
				8'h9C: decmult_11 = 8'h33;
				8'h9D: decmult_11 = 8'h38;
				8'h9E: decmult_11 = 8'h25;
				8'h9F: decmult_11 = 8'h2E;
				8'hA0: decmult_11 = 8'h8C;
				8'hA1: decmult_11 = 8'h87;
				8'hA2: decmult_11 = 8'h9A;
				8'hA3: decmult_11 = 8'h91;
				8'hA4: decmult_11 = 8'hA0;
				8'hA5: decmult_11 = 8'hAB;
				8'hA6: decmult_11 = 8'hB6;
				8'hA7: decmult_11 = 8'hBD;
				8'hA8: decmult_11 = 8'hD4;
				8'hA9: decmult_11 = 8'hDF;
				8'hAA: decmult_11 = 8'hC2;
				8'hAB: decmult_11 = 8'hC9;
				8'hAC: decmult_11 = 8'hF8;
				8'hAD: decmult_11 = 8'hF3;
				8'hAE: decmult_11 = 8'hEE;
				8'hAF: decmult_11 = 8'hE5;
				8'hB0: decmult_11 = 8'h3C;
				8'hB1: decmult_11 = 8'h37;
				8'hB2: decmult_11 = 8'h2A;
				8'hB3: decmult_11 = 8'h21;
				8'hB4: decmult_11 = 8'h10;
				8'hB5: decmult_11 = 8'h1B;
				8'hB6: decmult_11 = 8'h06;
				8'hB7: decmult_11 = 8'h0D;
				8'hB8: decmult_11 = 8'h64;
				8'hB9: decmult_11 = 8'h6F;
				8'hBA: decmult_11 = 8'h72;
				8'hBB: decmult_11 = 8'h79;
				8'hBC: decmult_11 = 8'h48;
				8'hBD: decmult_11 = 8'h43;
				8'hBE: decmult_11 = 8'h5E;
				8'hBF: decmult_11 = 8'h55;
				8'hC0: decmult_11 = 8'h01;
				8'hC1: decmult_11 = 8'h0A;
				8'hC2: decmult_11 = 8'h17;
				8'hC3: decmult_11 = 8'h1C;
				8'hC4: decmult_11 = 8'h2D;
				8'hC5: decmult_11 = 8'h26;
				8'hC6: decmult_11 = 8'h3B;
				8'hC7: decmult_11 = 8'h30;
				8'hC8: decmult_11 = 8'h59;
				8'hC9: decmult_11 = 8'h52;
				8'hCA: decmult_11 = 8'h4F;
				8'hCB: decmult_11 = 8'h44;
				8'hCC: decmult_11 = 8'h75;
				8'hCD: decmult_11 = 8'h7E;
				8'hCE: decmult_11 = 8'h63;
				8'hCF: decmult_11 = 8'h68;
				8'hD0: decmult_11 = 8'hB1;
				8'hD1: decmult_11 = 8'hBA;
				8'hD2: decmult_11 = 8'hA7;
				8'hD3: decmult_11 = 8'hAC;
				8'hD4: decmult_11 = 8'h9D;
				8'hD5: decmult_11 = 8'h96;
				8'hD6: decmult_11 = 8'h8B;
				8'hD7: decmult_11 = 8'h80;
				8'hD8: decmult_11 = 8'hE9;
				8'hD9: decmult_11 = 8'hE2;
				8'hDA: decmult_11 = 8'hFF;
				8'hDB: decmult_11 = 8'hF4;
				8'hDC: decmult_11 = 8'hC5;
				8'hDD: decmult_11 = 8'hCE;
				8'hDE: decmult_11 = 8'hD3;
				8'hDF: decmult_11 = 8'hD8;
				8'hE0: decmult_11 = 8'h7A;
				8'hE1: decmult_11 = 8'h71;
				8'hE2: decmult_11 = 8'h6C;
				8'hE3: decmult_11 = 8'h67;
				8'hE4: decmult_11 = 8'h56;
				8'hE5: decmult_11 = 8'h5D;
				8'hE6: decmult_11 = 8'h40;
				8'hE7: decmult_11 = 8'h4B;
				8'hE8: decmult_11 = 8'h22;
				8'hE9: decmult_11 = 8'h29;
				8'hEA: decmult_11 = 8'h34;
				8'hEB: decmult_11 = 8'h3F;
				8'hEC: decmult_11 = 8'h0E;
				8'hED: decmult_11 = 8'h05;
				8'hEE: decmult_11 = 8'h18;
				8'hEF: decmult_11 = 8'h13;
				8'hF0: decmult_11 = 8'hCA;
				8'hF1: decmult_11 = 8'hC1;
				8'hF2: decmult_11 = 8'hDC;
				8'hF3: decmult_11 = 8'hD7;
				8'hF4: decmult_11 = 8'hE6;
				8'hF5: decmult_11 = 8'hED;
				8'hF6: decmult_11 = 8'hF0;
				8'hF7: decmult_11 = 8'hFB;
				8'hF8: decmult_11 = 8'h92;
				8'hF9: decmult_11 = 8'h99;
				8'hFA: decmult_11 = 8'h84;
				8'hFB: decmult_11 = 8'h8F;
				8'hFC: decmult_11 = 8'hBE;
				8'hFD: decmult_11 = 8'hB5;
				8'hFE: decmult_11 = 8'hA8;
				8'hFF: decmult_11 = 8'hA3;
		  endcase
	 endfunction
	 
	 //function holding case statement multiply by 13
	 function [7:0] decmult_13(input [7:0] num);
		  case (num)
				8'h00: decmult_13 = 8'h00;
				8'h01: decmult_13 = 8'h0D;
				8'h02: decmult_13 = 8'h1A;
				8'h03: decmult_13 = 8'h17;
				8'h04: decmult_13 = 8'h34;
				8'h05: decmult_13 = 8'h39;
				8'h06: decmult_13 = 8'h2E;
				8'h07: decmult_13 = 8'h23;
				8'h08: decmult_13 = 8'h68;
				8'h09: decmult_13 = 8'h65;
				8'h0A: decmult_13 = 8'h72;
				8'h0B: decmult_13 = 8'h7F;
				8'h0C: decmult_13 = 8'h5C;
				8'h0D: decmult_13 = 8'h51;
				8'h0E: decmult_13 = 8'h46;
				8'h0F: decmult_13 = 8'h4B;
				8'h10: decmult_13 = 8'hD0;
				8'h11: decmult_13 = 8'hDD;
				8'h12: decmult_13 = 8'hCA;
				8'h13: decmult_13 = 8'hC7;
				8'h14: decmult_13 = 8'hE4;
				8'h15: decmult_13 = 8'hE9;
				8'h16: decmult_13 = 8'hFE;
				8'h17: decmult_13 = 8'hF3;
				8'h18: decmult_13 = 8'hB8;
				8'h19: decmult_13 = 8'hB5;
				8'h1A: decmult_13 = 8'hA2;
				8'h1B: decmult_13 = 8'hAF;
				8'h1C: decmult_13 = 8'h8C;
				8'h1D: decmult_13 = 8'h81;
				8'h1E: decmult_13 = 8'h96;
				8'h1F: decmult_13 = 8'h9B;
				8'h20: decmult_13 = 8'hBB;
				8'h21: decmult_13 = 8'hB6;
				8'h22: decmult_13 = 8'hA1;
				8'h23: decmult_13 = 8'hAC;
				8'h24: decmult_13 = 8'h8F;
				8'h25: decmult_13 = 8'h82;
				8'h26: decmult_13 = 8'h95;
				8'h27: decmult_13 = 8'h98;
				8'h28: decmult_13 = 8'hD3;
				8'h29: decmult_13 = 8'hDE;
				8'h2A: decmult_13 = 8'hC9;
				8'h2B: decmult_13 = 8'hC4;
				8'h2C: decmult_13 = 8'hE7;
				8'h2D: decmult_13 = 8'hEA;
				8'h2E: decmult_13 = 8'hFD;
				8'h2F: decmult_13 = 8'hF0;
				8'h30: decmult_13 = 8'h6B;
				8'h31: decmult_13 = 8'h66;
				8'h32: decmult_13 = 8'h71;
				8'h33: decmult_13 = 8'h7C;
				8'h34: decmult_13 = 8'h5F;
				8'h35: decmult_13 = 8'h52;
				8'h36: decmult_13 = 8'h45;
				8'h37: decmult_13 = 8'h48;
				8'h38: decmult_13 = 8'h03;
				8'h39: decmult_13 = 8'h0E;
				8'h3A: decmult_13 = 8'h19;
				8'h3B: decmult_13 = 8'h14;
				8'h3C: decmult_13 = 8'h37;
				8'h3D: decmult_13 = 8'h3A;
				8'h3E: decmult_13 = 8'h2D;
				8'h3F: decmult_13 = 8'h20;
				8'h40: decmult_13 = 8'h6D;
				8'h41: decmult_13 = 8'h60;
				8'h42: decmult_13 = 8'h77;
				8'h43: decmult_13 = 8'h7A;
				8'h44: decmult_13 = 8'h59;
				8'h45: decmult_13 = 8'h54;
				8'h46: decmult_13 = 8'h43;
				8'h47: decmult_13 = 8'h4E;
				8'h48: decmult_13 = 8'h05;
				8'h49: decmult_13 = 8'h08;
				8'h4A: decmult_13 = 8'h1F;
				8'h4B: decmult_13 = 8'h12;
				8'h4C: decmult_13 = 8'h31;
				8'h4D: decmult_13 = 8'h3C;
				8'h4E: decmult_13 = 8'h2B;
				8'h4F: decmult_13 = 8'h26;
				8'h50: decmult_13 = 8'hBD;
				8'h51: decmult_13 = 8'hB0;
				8'h52: decmult_13 = 8'hA7;
				8'h53: decmult_13 = 8'hAA;
				8'h54: decmult_13 = 8'h89;
				8'h55: decmult_13 = 8'h84;
				8'h56: decmult_13 = 8'h93;
				8'h57: decmult_13 = 8'h9E;
				8'h58: decmult_13 = 8'hD5;
				8'h59: decmult_13 = 8'hD8;
				8'h5A: decmult_13 = 8'hCF;
				8'h5B: decmult_13 = 8'hC2;
				8'h5C: decmult_13 = 8'hE1;
				8'h5D: decmult_13 = 8'hEC;
				8'h5E: decmult_13 = 8'hFB;
				8'h5F: decmult_13 = 8'hF6;
				8'h60: decmult_13 = 8'hD6;
				8'h61: decmult_13 = 8'hDB;
				8'h62: decmult_13 = 8'hCC;
				8'h63: decmult_13 = 8'hC1;
				8'h64: decmult_13 = 8'hE2;
				8'h65: decmult_13 = 8'hEF;
				8'h66: decmult_13 = 8'hF8;
				8'h67: decmult_13 = 8'hF5;
				8'h68: decmult_13 = 8'hBE;
				8'h69: decmult_13 = 8'hB3;
				8'h6A: decmult_13 = 8'hA4;
				8'h6B: decmult_13 = 8'hA9;
				8'h6C: decmult_13 = 8'h8A;
				8'h6D: decmult_13 = 8'h87;
				8'h6E: decmult_13 = 8'h90;
				8'h6F: decmult_13 = 8'h9D;
				8'h70: decmult_13 = 8'h06;
				8'h71: decmult_13 = 8'h0B;
				8'h72: decmult_13 = 8'h1C;
				8'h73: decmult_13 = 8'h11;
				8'h74: decmult_13 = 8'h32;
				8'h75: decmult_13 = 8'h3F;
				8'h76: decmult_13 = 8'h28;
				8'h77: decmult_13 = 8'h25;
				8'h78: decmult_13 = 8'h6E;
				8'h79: decmult_13 = 8'h63;
				8'h7A: decmult_13 = 8'h74;
				8'h7B: decmult_13 = 8'h79;
				8'h7C: decmult_13 = 8'h5A;
				8'h7D: decmult_13 = 8'h57;
				8'h7E: decmult_13 = 8'h40;
				8'h7F: decmult_13 = 8'h4D;
				8'h80: decmult_13 = 8'hDA;
				8'h81: decmult_13 = 8'hD7;
				8'h82: decmult_13 = 8'hC0;
				8'h83: decmult_13 = 8'hCD;
				8'h84: decmult_13 = 8'hEE;
				8'h85: decmult_13 = 8'hE3;
				8'h86: decmult_13 = 8'hF4;
				8'h87: decmult_13 = 8'hF9;
				8'h88: decmult_13 = 8'hB2;
				8'h89: decmult_13 = 8'hBF;
				8'h8A: decmult_13 = 8'hA8;
				8'h8B: decmult_13 = 8'hA5;
				8'h8C: decmult_13 = 8'h86;
				8'h8D: decmult_13 = 8'h8B;
				8'h8E: decmult_13 = 8'h9C;
				8'h8F: decmult_13 = 8'h91;
				8'h90: decmult_13 = 8'h0A;
				8'h91: decmult_13 = 8'h07;
				8'h92: decmult_13 = 8'h10;
				8'h93: decmult_13 = 8'h1D;
				8'h94: decmult_13 = 8'h3E;
				8'h95: decmult_13 = 8'h33;
				8'h96: decmult_13 = 8'h24;
				8'h97: decmult_13 = 8'h29;
				8'h98: decmult_13 = 8'h62;
				8'h99: decmult_13 = 8'h6F;
				8'h9A: decmult_13 = 8'h78;
				8'h9B: decmult_13 = 8'h75;
				8'h9C: decmult_13 = 8'h56;
				8'h9D: decmult_13 = 8'h5B;
				8'h9E: decmult_13 = 8'h4C;
				8'h9F: decmult_13 = 8'h41;
				8'hA0: decmult_13 = 8'h61;
				8'hA1: decmult_13 = 8'h6C;
				8'hA2: decmult_13 = 8'h7B;
				8'hA3: decmult_13 = 8'h76;
				8'hA4: decmult_13 = 8'h55;
				8'hA5: decmult_13 = 8'h58;
				8'hA6: decmult_13 = 8'h4F;
				8'hA7: decmult_13 = 8'h42;
				8'hA8: decmult_13 = 8'h09;
				8'hA9: decmult_13 = 8'h04;
				8'hAA: decmult_13 = 8'h13;
				8'hAB: decmult_13 = 8'h1E;
				8'hAC: decmult_13 = 8'h3D;
				8'hAD: decmult_13 = 8'h30;
				8'hAE: decmult_13 = 8'h27;
				8'hAF: decmult_13 = 8'h2A;
				8'hB0: decmult_13 = 8'hB1;
				8'hB1: decmult_13 = 8'hBC;
				8'hB2: decmult_13 = 8'hAB;
				8'hB3: decmult_13 = 8'hA6;
				8'hB4: decmult_13 = 8'h85;
				8'hB5: decmult_13 = 8'h88;
				8'hB6: decmult_13 = 8'h9F;
				8'hB7: decmult_13 = 8'h92;
				8'hB8: decmult_13 = 8'hD9;
				8'hB9: decmult_13 = 8'hD4;
				8'hBA: decmult_13 = 8'hC3;
				8'hBB: decmult_13 = 8'hCE;
				8'hBC: decmult_13 = 8'hED;
				8'hBD: decmult_13 = 8'hE0;
				8'hBE: decmult_13 = 8'hF7;
				8'hBF: decmult_13 = 8'hFA;
				8'hC0: decmult_13 = 8'hB7;
				8'hC1: decmult_13 = 8'hBA;
				8'hC2: decmult_13 = 8'hAD;
				8'hC3: decmult_13 = 8'hA0;
				8'hC4: decmult_13 = 8'h83;
				8'hC5: decmult_13 = 8'h8E;
				8'hC6: decmult_13 = 8'h99;
				8'hC7: decmult_13 = 8'h94;
				8'hC8: decmult_13 = 8'hDF;
				8'hC9: decmult_13 = 8'hD2;
				8'hCA: decmult_13 = 8'hC5;
				8'hCB: decmult_13 = 8'hC8;
				8'hCC: decmult_13 = 8'hEB;
				8'hCD: decmult_13 = 8'hE6;
				8'hCE: decmult_13 = 8'hF1;
				8'hCF: decmult_13 = 8'hFC;
				8'hD0: decmult_13 = 8'h67;
				8'hD1: decmult_13 = 8'h6A;
				8'hD2: decmult_13 = 8'h7D;
				8'hD3: decmult_13 = 8'h70;
				8'hD4: decmult_13 = 8'h53;
				8'hD5: decmult_13 = 8'h5E;
				8'hD6: decmult_13 = 8'h49;
				8'hD7: decmult_13 = 8'h44;
				8'hD8: decmult_13 = 8'h0F;
				8'hD9: decmult_13 = 8'h02;
				8'hDA: decmult_13 = 8'h15;
				8'hDB: decmult_13 = 8'h18;
				8'hDC: decmult_13 = 8'h3B;
				8'hDD: decmult_13 = 8'h36;
				8'hDE: decmult_13 = 8'h21;
				8'hDF: decmult_13 = 8'h2C;
				8'hE0: decmult_13 = 8'h0C;
				8'hE1: decmult_13 = 8'h01;
				8'hE2: decmult_13 = 8'h16;
				8'hE3: decmult_13 = 8'h1B;
				8'hE4: decmult_13 = 8'h38;
				8'hE5: decmult_13 = 8'h35;
				8'hE6: decmult_13 = 8'h22;
				8'hE7: decmult_13 = 8'h2F;
				8'hE8: decmult_13 = 8'h64;
				8'hE9: decmult_13 = 8'h69;
				8'hEA: decmult_13 = 8'h7E;
				8'hEB: decmult_13 = 8'h73;
				8'hEC: decmult_13 = 8'h50;
				8'hED: decmult_13 = 8'h5D;
				8'hEE: decmult_13 = 8'h4A;
				8'hEF: decmult_13 = 8'h47;
				8'hF0: decmult_13 = 8'hDC;
				8'hF1: decmult_13 = 8'hD1;
				8'hF2: decmult_13 = 8'hC6;
				8'hF3: decmult_13 = 8'hCB;
				8'hF4: decmult_13 = 8'hE8;
				8'hF5: decmult_13 = 8'hE5;
				8'hF6: decmult_13 = 8'hF2;
				8'hF7: decmult_13 = 8'hFF;
				8'hF8: decmult_13 = 8'hB4;
				8'hF9: decmult_13 = 8'hB9;
				8'hFA: decmult_13 = 8'hAE;
				8'hFB: decmult_13 = 8'hA3;
				8'hFC: decmult_13 = 8'h80;
				8'hFD: decmult_13 = 8'h8D;
				8'hFE: decmult_13 = 8'h9A;
				8'hFF: decmult_13 = 8'h97;
		  endcase
	 endfunction
	 
	 //function holding case statement multiply by 14
	 function [7:0] decmult_14(input [7:0] num);
		  case (num)
				8'h00: decmult_14 = 8'h00;
				8'h01: decmult_14 = 8'h0E;
				8'h02: decmult_14 = 8'h1C;
				8'h03: decmult_14 = 8'h12;
				8'h04: decmult_14 = 8'h38;
				8'h05: decmult_14 = 8'h36;
				8'h06: decmult_14 = 8'h24;
				8'h07: decmult_14 = 8'h2A;
				8'h08: decmult_14 = 8'h70;
				8'h09: decmult_14 = 8'h7E;
				8'h0A: decmult_14 = 8'h6C;
				8'h0B: decmult_14 = 8'h62;
				8'h0C: decmult_14 = 8'h48;
				8'h0D: decmult_14 = 8'h46;
				8'h0E: decmult_14 = 8'h54;
				8'h0F: decmult_14 = 8'h5A;
				8'h10: decmult_14 = 8'hE0;
				8'h11: decmult_14 = 8'hEE;
				8'h12: decmult_14 = 8'hFC;
				8'h13: decmult_14 = 8'hF2;
				8'h14: decmult_14 = 8'hD8;
				8'h15: decmult_14 = 8'hD6;
				8'h16: decmult_14 = 8'hC4;
				8'h17: decmult_14 = 8'hCA;
				8'h18: decmult_14 = 8'h90;
				8'h19: decmult_14 = 8'h9E;
				8'h1A: decmult_14 = 8'h8C;
				8'h1B: decmult_14 = 8'h82;
				8'h1C: decmult_14 = 8'hA8;
				8'h1D: decmult_14 = 8'hA6;
				8'h1E: decmult_14 = 8'hB4;
				8'h1F: decmult_14 = 8'hBA;
				8'h20: decmult_14 = 8'hDB;
				8'h21: decmult_14 = 8'hD5;
				8'h22: decmult_14 = 8'hC7;
				8'h23: decmult_14 = 8'hC9;
				8'h24: decmult_14 = 8'hE3;
				8'h25: decmult_14 = 8'hED;
				8'h26: decmult_14 = 8'hFF;
				8'h27: decmult_14 = 8'hF1;
				8'h28: decmult_14 = 8'hAB;
				8'h29: decmult_14 = 8'hA5;
				8'h2A: decmult_14 = 8'hB7;
				8'h2B: decmult_14 = 8'hB9;
				8'h2C: decmult_14 = 8'h93;
				8'h2D: decmult_14 = 8'h9D;
				8'h2E: decmult_14 = 8'h8F;
				8'h2F: decmult_14 = 8'h81;
				8'h30: decmult_14 = 8'h3B;
				8'h31: decmult_14 = 8'h35;
				8'h32: decmult_14 = 8'h27;
				8'h33: decmult_14 = 8'h29;
				8'h34: decmult_14 = 8'h03;
				8'h35: decmult_14 = 8'h0D;
				8'h36: decmult_14 = 8'h1F;
				8'h37: decmult_14 = 8'h11;
				8'h38: decmult_14 = 8'h4B;
				8'h39: decmult_14 = 8'h45;
				8'h3A: decmult_14 = 8'h57;
				8'h3B: decmult_14 = 8'h59;
				8'h3C: decmult_14 = 8'h73;
				8'h3D: decmult_14 = 8'h7D;
				8'h3E: decmult_14 = 8'h6F;
				8'h3F: decmult_14 = 8'h61;
				8'h40: decmult_14 = 8'hAD;
				8'h41: decmult_14 = 8'hA3;
				8'h42: decmult_14 = 8'hB1;
				8'h43: decmult_14 = 8'hBF;
				8'h44: decmult_14 = 8'h95;
				8'h45: decmult_14 = 8'h9B;
				8'h46: decmult_14 = 8'h89;
				8'h47: decmult_14 = 8'h87;
				8'h48: decmult_14 = 8'hDD;
				8'h49: decmult_14 = 8'hD3;
				8'h4A: decmult_14 = 8'hC1;
				8'h4B: decmult_14 = 8'hCF;
				8'h4C: decmult_14 = 8'hE5;
				8'h4D: decmult_14 = 8'hEB;
				8'h4E: decmult_14 = 8'hF9;
				8'h4F: decmult_14 = 8'hF7;
				8'h50: decmult_14 = 8'h4D;
				8'h51: decmult_14 = 8'h43;
				8'h52: decmult_14 = 8'h51;
				8'h53: decmult_14 = 8'h5F;
				8'h54: decmult_14 = 8'h75;
				8'h55: decmult_14 = 8'h7B;
				8'h56: decmult_14 = 8'h69;
				8'h57: decmult_14 = 8'h67;
				8'h58: decmult_14 = 8'h3D;
				8'h59: decmult_14 = 8'h33;
				8'h5A: decmult_14 = 8'h21;
				8'h5B: decmult_14 = 8'h2F;
				8'h5C: decmult_14 = 8'h05;
				8'h5D: decmult_14 = 8'h0B;
				8'h5E: decmult_14 = 8'h19;
				8'h5F: decmult_14 = 8'h17;
				8'h60: decmult_14 = 8'h76;
				8'h61: decmult_14 = 8'h78;
				8'h62: decmult_14 = 8'h6A;
				8'h63: decmult_14 = 8'h64;
				8'h64: decmult_14 = 8'h4E;
				8'h65: decmult_14 = 8'h40;
				8'h66: decmult_14 = 8'h52;
				8'h67: decmult_14 = 8'h5C;
				8'h68: decmult_14 = 8'h06;
				8'h69: decmult_14 = 8'h08;
				8'h6A: decmult_14 = 8'h1A;
				8'h6B: decmult_14 = 8'h14;
				8'h6C: decmult_14 = 8'h3E;
				8'h6D: decmult_14 = 8'h30;
				8'h6E: decmult_14 = 8'h22;
				8'h6F: decmult_14 = 8'h2C;
				8'h70: decmult_14 = 8'h96;
				8'h71: decmult_14 = 8'h98;
				8'h72: decmult_14 = 8'h8A;
				8'h73: decmult_14 = 8'h84;
				8'h74: decmult_14 = 8'hAE;
				8'h75: decmult_14 = 8'hA0;
				8'h76: decmult_14 = 8'hB2;
				8'h77: decmult_14 = 8'hBC;
				8'h78: decmult_14 = 8'hE6;
				8'h79: decmult_14 = 8'hE8;
				8'h7A: decmult_14 = 8'hFA;
				8'h7B: decmult_14 = 8'hF4;
				8'h7C: decmult_14 = 8'hDE;
				8'h7D: decmult_14 = 8'hD0;
				8'h7E: decmult_14 = 8'hC2;
				8'h7F: decmult_14 = 8'hCC;
				8'h80: decmult_14 = 8'h41;
				8'h81: decmult_14 = 8'h4F;
				8'h82: decmult_14 = 8'h5D;
				8'h83: decmult_14 = 8'h53;
				8'h84: decmult_14 = 8'h79;
				8'h85: decmult_14 = 8'h77;
				8'h86: decmult_14 = 8'h65;
				8'h87: decmult_14 = 8'h6B;
				8'h88: decmult_14 = 8'h31;
				8'h89: decmult_14 = 8'h3F;
				8'h8A: decmult_14 = 8'h2D;
				8'h8B: decmult_14 = 8'h23;
				8'h8C: decmult_14 = 8'h09;
				8'h8D: decmult_14 = 8'h07;
				8'h8E: decmult_14 = 8'h15;
				8'h8F: decmult_14 = 8'h1B;
				8'h90: decmult_14 = 8'hA1;
				8'h91: decmult_14 = 8'hAF;
				8'h92: decmult_14 = 8'hBD;
				8'h93: decmult_14 = 8'hB3;
				8'h94: decmult_14 = 8'h99;
				8'h95: decmult_14 = 8'h97;
				8'h96: decmult_14 = 8'h85;
				8'h97: decmult_14 = 8'h8B;
				8'h98: decmult_14 = 8'hD1;
				8'h99: decmult_14 = 8'hDF;
				8'h9A: decmult_14 = 8'hCD;
				8'h9B: decmult_14 = 8'hC3;
				8'h9C: decmult_14 = 8'hE9;
				8'h9D: decmult_14 = 8'hE7;
				8'h9E: decmult_14 = 8'hF5;
				8'h9F: decmult_14 = 8'hFB;
				8'hA0: decmult_14 = 8'h9A;
				8'hA1: decmult_14 = 8'h94;
				8'hA2: decmult_14 = 8'h86;
				8'hA3: decmult_14 = 8'h88;
				8'hA4: decmult_14 = 8'hA2;
				8'hA5: decmult_14 = 8'hAC;
				8'hA6: decmult_14 = 8'hBE;
				8'hA7: decmult_14 = 8'hB0;
				8'hA8: decmult_14 = 8'hEA;
				8'hA9: decmult_14 = 8'hE4;
				8'hAA: decmult_14 = 8'hF6;
				8'hAB: decmult_14 = 8'hF8;
				8'hAC: decmult_14 = 8'hD2;
				8'hAD: decmult_14 = 8'hDC;
				8'hAE: decmult_14 = 8'hCE;
				8'hAF: decmult_14 = 8'hC0;
				8'hB0: decmult_14 = 8'h7A;
				8'hB1: decmult_14 = 8'h74;
				8'hB2: decmult_14 = 8'h66;
				8'hB3: decmult_14 = 8'h68;
				8'hB4: decmult_14 = 8'h42;
				8'hB5: decmult_14 = 8'h4C;
				8'hB6: decmult_14 = 8'h5E;
				8'hB7: decmult_14 = 8'h50;
				8'hB8: decmult_14 = 8'h0A;
				8'hB9: decmult_14 = 8'h04;
				8'hBA: decmult_14 = 8'h16;
				8'hBB: decmult_14 = 8'h18;
				8'hBC: decmult_14 = 8'h32;
				8'hBD: decmult_14 = 8'h3C;
				8'hBE: decmult_14 = 8'h2E;
				8'hBF: decmult_14 = 8'h20;
				8'hC0: decmult_14 = 8'hEC;
				8'hC1: decmult_14 = 8'hE2;
				8'hC2: decmult_14 = 8'hF0;
				8'hC3: decmult_14 = 8'hFE;
				8'hC4: decmult_14 = 8'hD4;
				8'hC5: decmult_14 = 8'hDA;
				8'hC6: decmult_14 = 8'hC8;
				8'hC7: decmult_14 = 8'hC6;
				8'hC8: decmult_14 = 8'h9C;
				8'hC9: decmult_14 = 8'h92;
				8'hCA: decmult_14 = 8'h80;
				8'hCB: decmult_14 = 8'h8E;
				8'hCC: decmult_14 = 8'hA4;
				8'hCD: decmult_14 = 8'hAA;
				8'hCE: decmult_14 = 8'hB8;
				8'hCF: decmult_14 = 8'hB6;
				8'hD0: decmult_14 = 8'h0C;
				8'hD1: decmult_14 = 8'h02;
				8'hD2: decmult_14 = 8'h10;
				8'hD3: decmult_14 = 8'h1E;
				8'hD4: decmult_14 = 8'h34;
				8'hD5: decmult_14 = 8'h3A;
				8'hD6: decmult_14 = 8'h28;
				8'hD7: decmult_14 = 8'h26;
				8'hD8: decmult_14 = 8'h7C;
				8'hD9: decmult_14 = 8'h72;
				8'hDA: decmult_14 = 8'h60;
				8'hDB: decmult_14 = 8'h6E;
				8'hDC: decmult_14 = 8'h44;
				8'hDD: decmult_14 = 8'h4A;
				8'hDE: decmult_14 = 8'h58;
				8'hDF: decmult_14 = 8'h56;
				8'hE0: decmult_14 = 8'h37;
				8'hE1: decmult_14 = 8'h39;
				8'hE2: decmult_14 = 8'h2B;
				8'hE3: decmult_14 = 8'h25;
				8'hE4: decmult_14 = 8'h0F;
				8'hE5: decmult_14 = 8'h01;
				8'hE6: decmult_14 = 8'h13;
				8'hE7: decmult_14 = 8'h1D;
				8'hE8: decmult_14 = 8'h47;
				8'hE9: decmult_14 = 8'h49;
				8'hEA: decmult_14 = 8'h5B;
				8'hEB: decmult_14 = 8'h55;
				8'hEC: decmult_14 = 8'h7F;
				8'hED: decmult_14 = 8'h71;
				8'hEE: decmult_14 = 8'h63;
				8'hEF: decmult_14 = 8'h6D;
				8'hF0: decmult_14 = 8'hD7;
				8'hF1: decmult_14 = 8'hD9;
				8'hF2: decmult_14 = 8'hCB;
				8'hF3: decmult_14 = 8'hC5;
				8'hF4: decmult_14 = 8'hEF;
				8'hF5: decmult_14 = 8'hE1;
				8'hF6: decmult_14 = 8'hF3;
				8'hF7: decmult_14 = 8'hFD;
				8'hF8: decmult_14 = 8'hA7;
				8'hF9: decmult_14 = 8'hA9;
				8'hFA: decmult_14 = 8'hBB;
				8'hFB: decmult_14 = 8'hB5;
				8'hFC: decmult_14 = 8'h9F;
				8'hFD: decmult_14 = 8'h91;
				8'hFE: decmult_14 = 8'h83;
				8'hFF: decmult_14 = 8'h8D;
		  endcase
	 endfunction
endmodule
